module  lab8 		( input         CLOCK_50,
                       input[3:0]    KEY, //bit 0 is set up as Reset
							  output [6:0]  HEX0, HEX1, HEX6, HEX7,HEX5,HEX4,
							  //output [8:0]  LEDG,
							  //output [17:0] LEDR,
							  // VGA Interface 
                       output [7:0]  VGA_R,					//VGA Red
							                VGA_G,					//VGA Green
												 VGA_B,					//VGA Blue
							  output        VGA_CLK,				//VGA Clock
							                VGA_SYNC_N,			//VGA Sync signal
												 VGA_BLANK_N,			//VGA Blank signal
												 VGA_VS,					//VGA virtical sync signal	
												 VGA_HS,					//VGA horizontal sync signal
							  // CY7C67200 Interface
							  inout [15:0]  OTG_DATA,						//	CY7C67200 Data bus 16 Bits
							  output [1:0]  OTG_ADDR,						//	CY7C67200 Address 2 Bits
							  output        OTG_CS_N,						//	CY7C67200 Chip Select
												 OTG_RD_N,						//	CY7C67200 Write
												 OTG_WR_N,						//	CY7C67200 Read
												 OTG_RST_N,						//	CY7C67200 Reset
							  input			 OTG_INT,						//	CY7C67200 Interrupt
							  // SDRAM Interface for Nios II Software
							  output [12:0] DRAM_ADDR,				// SDRAM Address 13 Bits
							  inout [31:0]  DRAM_DQ,				// SDRAM Data 32 Bits
							  output [1:0]  DRAM_BA,				// SDRAM Bank Address 2 Bits
							  output [3:0]  DRAM_DQM,				// SDRAM Data Mast 4 Bits
							  output			 DRAM_RAS_N,			// SDRAM Row Address Strobe
							  output			 DRAM_CAS_N,			// SDRAM Column Address Strobe
							  output			 DRAM_CKE,				// SDRAM Clock Enable
							  output			 DRAM_WE_N,				// SDRAM Write Enable
							  output			 DRAM_CS_N,				// SDRAM Chip Select
							  output			 DRAM_CLK				// SDRAM Clock
											);
    
    	logic Reset_h, vssig, Clk;
    	logic [9:0] drawxsig, drawysig, ballxsig, ballysig, ballsizesig, jumpxsig, jumpysig, jumpsizesig, puckx, pucky, pucksize, WallballS, WallballX, WallballY;
		logic [15:0] keycode;
		logic MainS, StartScreen, Instructions, PauseScreen1, PauseScreen2, Game1Screen, Game2Screen, ExitScreen, Ready, Hoop;
		logic hit_floor, hit_target;
		logic [0:95][0:172][0:1] Title;
		logic [0:53][0:205][0:1] Names;
		logic [0:95][0:137][0:1] InstructionTXT;
		logic [0:25][0:116][0:1] MainOptions;
		logic [0:25][0:98][0:1] GameSelect;
		logic [0:150][0:126][0:3] HoopTXT;
		logic [0:47][0:63][0:1] PauseTXT;
		logic [0:399][0:9][0:1] wallTXT;


		logic [10:0] Score;
		logic [3:0] hextotal, hextotal2, hextotal3, hextotal4;   



	assign Clk = CLOCK_50;
    	assign {Reset_h}=~ (KEY[0]);  // The push buttons are active low
	
	wire [1:0] hpi_addr;
	wire [15:0] hpi_data_in, hpi_data_out;
	wire hpi_r, hpi_w,hpi_cs;
	 


	 hpi_io_intf hpi_io_inst(   .from_sw_address(hpi_addr),
										 .from_sw_data_in(hpi_data_in),
										 .from_sw_data_out(hpi_data_out),
										 .from_sw_r(hpi_r),
										 .from_sw_w(hpi_w),
										 .from_sw_cs(hpi_cs),
		 								 .OTG_DATA(OTG_DATA),    
										 .OTG_ADDR(OTG_ADDR),    
										 .OTG_RD_N(OTG_RD_N),    
										 .OTG_WR_N(OTG_WR_N),    
										 .OTG_CS_N(OTG_CS_N),    
										 .OTG_RST_N(OTG_RST_N),   
										 .OTG_INT(OTG_INT),
										 .Clk(Clk),
										 .Reset(Reset_h)
	 );
	 
	 //The connections for nios_system might be named different depending on how you set up Qsys
	 lab8_soc nios_system(
										 .clk_clk(Clk),         
										 .reset_reset_n(KEY[0]),   
										 .sdram_wire_addr(DRAM_ADDR), 
										 .sdram_wire_ba(DRAM_BA),   
										 .sdram_wire_cas_n(DRAM_CAS_N),
										 .sdram_wire_cke(DRAM_CKE),  
										 .sdram_wire_cs_n(DRAM_CS_N), 
										 .sdram_wire_dq(DRAM_DQ),   
										 .sdram_wire_dqm(DRAM_DQM),  
										 .sdram_wire_ras_n(DRAM_RAS_N),
										 .sdram_wire_we_n(DRAM_WE_N), 
										 .sdram_clk_clk(DRAM_CLK),
										 .keycode_export(keycode),  
										 .otg_hpi_address_export(hpi_addr),
										 .otg_hpi_data_in_port(hpi_data_in),
										 .otg_hpi_data_out_port(hpi_data_out),
										 .otg_hpi_cs_export(hpi_cs),
										 .otg_hpi_r_export(hpi_r),
										 .otg_hpi_w_export(hpi_w));
										 
	//Fill in the connections for the rest of the modules 
  	vga_controller vgasync_instance( .Clk(Clk),
												.Reset(Reset_h),
												.hs(VGA_HS),
												.vs(VGA_VS),
												.pixel_clk(VGA_CLK),
												.blank(VGA_BLANK_N),
												.sync(VGA_SYNC_N),
												.DrawX(drawxsig),
												.DrawY(drawysig)
					);
							
   slime1 player1( .Reset(Reset_h),
								.frame_clk(VGA_VS),
								.key(keycode),
								.BallX(ballxsig),
								.BallY(ballysig),
								.BallS(ballsizesig)
					);
								
	slime2 player2( .Reset(Reset_h),
								.frame_clk(VGA_VS),
								.key1(!KEY[1]),
								.key2(!KEY[2]),
								.key3(!KEY[3]),
								.JumpX(jumpxsig),
								.JumpY(jumpysig),
								.JumpS(jumpsizesig)
					);
										
	puck  puckinstance (
								.Reset(Reset_h), 
								.frame_clk(VGA_VS),
								.Actor_X(ballxsig), 
								.Actor_Y(ballysig), 
								.Actor_Size(ballsizesig), 
								.Jump_X(jumpxsig), 
								.Jump_Y(jumpysig), 
								.Jump_Size(jumpsizesig),
								.BallX(puckx), 
								.BallY(pucky), 
								.BallS(pucksize),
								.hit_floor(hit_floor), 
								.hit_target(hit_target),
								.hextotal(hextotal),
								.hextotal2(hextotal2),
								.Game1Screen(Game1Screen), 
								.Game2Screen(Game2Screen)
								);
								
	wallball  wallbinstance (
								.Reset(Reset_h), 
								.frame_clk(VGA_VS),
								.Actor_X(ballxsig), 
								.Actor_Y(ballysig), 
								.Actor_Size(ballsizesig), 
								.BallX(WallballX), 
								.BallY(WallballY), 
								.BallS(WallballS),
								.hit_floor(hit_floor), 
								.hit_target(hit_target),
								.hextotal(hextotal3),
								.hextotal2(hextotal4)					
								);	

	color_mapper color_instance(	.JumpX(jumpxsig),
					.JumpY(jumpysig),
					.JumpS(jumpsizesig),
					.BallX(ballxsig),
					.BallY(ballysig),
					.DrawX(drawxsig),
					.DrawY(drawysig),
					.Ball_size(ballsizesig),
					.PuckX(puckx),
					.PuckY(pucky),
					.PuckS(pucksize),
					.WallballX(WallballX),
					.WallballY(WallballY),
					.WallballS(WallballS),
					.Red(VGA_R),
					.Green(VGA_G),
					.Blue(VGA_B),
					.Hoop(HoopTXT),
					.MainS(MainS),
					.StartScreen(StartScreen),
					.Instructions(Instructions),
					.PauseScreen1(PauseScreen1),
					.PauseScreen2(PauseScreen2),
					.Game1Screen(Game1Screen),
					.Game2Screen(Game2Screen),
					.ExitScreen(ExitScreen),
					.Ready(Ready),
					.Title(Title),
					.Names(Names),
					.InstructionTXT(InstructionTXT),
					.MainOptions(MainOptions),
					.GameSelect(GameSelect),
					.Pause(PauseTXT)
					);
	 

	gamelogic logic_instance ( 	.Reset(Reset_h), 
					.frame_clk(VGA_VS),
					.key(keycode),
					.MainS(MainS),
					.StartScreen(StartScreen),
					.Instructions(Instructions),
					.PauseScreen1(PauseScreen1),
					.PauseScreen2(PauseScreen2),
					.Game1Screen(Game1Screen),
					.Game2Screen(Game2Screen),
					.ExitScreen(ExitScreen),
					.hit_floor(hit_floor), 
					.hextotal(),
					.hextotal2(),
					.hit_target(hit_target),
					.Score(Score)
					);
					
	sprite_table spriteinstance (	.clk(VGA_VS),
											.Title(Title),
											.Names(Names),
											.Instructions(InstructionTXT),
											.MainOptions(MainOptions),
											.GameSelect(GameSelect),
											.Hoop(HoopTXT),
											.Pause(PauseTXT),
											.wall(wallTXT)
										);



	HexDriver hex_inst_0 (keycode[3:0], HEX0);
	HexDriver hex_inst_1 (keycode[7:4], HEX1);							  
	HexDriver hex_inst_2 (hextotal, HEX6);
	HexDriver hex_inst_3 (hextotal2, HEX7);
	HexDriver hex_inst_4 (hextotal3, HEX4);
	HexDriver hex_inst_5 (hextotal4, HEX5);

endmodule
